library STD;
library IEEE;
use IEEE.std_logic_1164.all;

entity and3 is
  port (
    x  : in  std_logic;
    y   : in  std_logic;
    z   : in  std_logic;
    o  : out std_logic
  );
end and3;

architecture structural of and3 is

  -- base 2-input AND gate
  component and2
    port (
      input0   : in  std_logic;
      input1   : in  std_logic;
      output0  : out std_logic
    );
  end component;

  -- internal signal
  signal t1 : std_logic;

begin
  -- first stage
  and2_0 : and2 port map(input0 => x, input1 => y, output0 => t1);

  -- second stage
  and2_1 : and2 port map(input0 => t1, input1 => z, output0 => o);

end structural;

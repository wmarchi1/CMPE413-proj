--
-- Entity: and2
-- Architecture : structural
-- Author: cpatel2
-- Created On: 11/11/2003
--
library STD;
library IEEE;
use IEEE.std_logic_1164.all;

entity and2 is

  port (
    input0   : in  std_logic;
    input1   : in  std_logic;
    output0   : out std_logic);
end and2;

architecture structural of and2 is

begin

  output <= input2 and input1;

end structural;
